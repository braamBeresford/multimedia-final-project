module quantization(input  logic clk,
		    input  logic start,
                    input  logic [7:0][7:0][9:0] in_matrix,
	            output logic [7:0][7:0][9:0] out_matrix,
	    	    output logic done);

endmodule	
